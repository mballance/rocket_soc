/****************************************************************************
 * RocketBFMBinds.sv
 ****************************************************************************/

/**
 * Module: RocketBFMBinds
 * 
 * TODO: Add module documentation
 */
module RocketBFMBinds;



endmodule


