

`include "uvm_macros.svh"
package rocket_soc_tests_pkg;
	import uvm_pkg::*;
	import rocket_soc_env_pkg::*;
	import vmon_client_pkg::*;
	import vmon_client_uvm_pkg::*;
	import uart_serial_agent_pkg::*;
	
	`include "rocket_soc_test_base.svh"
	
endpackage
