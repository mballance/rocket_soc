
`include "uvm_macros.svh"

package rocket_soc_subsys_env_pkg;
	import uvm_pkg::*;
	import hella_cache_master_agent_pkg::*;

	`include "rocket_soc_subsys_env.svh"
	
endpackage
