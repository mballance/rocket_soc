/****************************************************************************
 * RocketSocEnvTBBasePkg.sv
 ****************************************************************************/
`include "uvm_macros.svh"
/**
 * Package: RocketSocEnvBasePkg
 * 
 * TODO: Add package documentation
 */
package RocketSocTBEnvBasePkg;
	import uvm_pkg::*;
	import uart_serial_agent_pkg::*;
	
	`include "RocketSocTBEnvBase.svh"


endpackage


