
`include "uvm_macros.svh"

package rocket_soc_subsys_env_pkg;
	import uvm_pkg::*;
	import hella_cache_master_agent_pkg::*;
	import sv_bfms_api_pkg::*;
	import uex_pkg::*;
	import uart_serial_agent_pkg::*;
	import event_agent_pkg::*;
	import vmon_client_pkg::*;
	import vmon_client_uvm_pkg::*;
	import vmon_client_api_pkg::*;
	import uvmdev_vmon_pkg::*;

	`include "rocket_soc_subsys_mem_services.svh"
	`include "rocket_soc_subsys_env.svh"
	
endpackage
