/****************************************************************************
 * rocket_soc_subsys_tb.sv
 ****************************************************************************/

/**
 * Module: rocket_soc_subsys_tb
 * 
 * TODO: Add module documentation
 */
`include "uvm_macros.svh"
module rocket_soc_subsys_tb;
	import uvm_pkg::*;
	import rocket_soc_subsys_tests_pkg::*;
	
	rocket_soc_tb tb();
	
//	initial begin
//		run_test();
//	end

endmodule

