
`include "uvm_macros.svh"

package rocket_soc_subsys_env_pkg;
	import uvm_pkg::*;
	import hella_cache_master_agent_pkg::*;
	import sv_bfms_api_pkg::*;
	import uex_pkg::*;

	`include "rocket_soc_subsys_mem_services.svh"
	`include "rocket_soc_subsys_env.svh"
	
endpackage
