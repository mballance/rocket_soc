

`include "uvm_macros.svh"
package rocket_soc_subsys_tests_pkg;
	import uvm_pkg::*;
	import rocket_soc_subsys_env_pkg::*;
	
	`include "rocket_soc_subsys_test_base.svh"
	
endpackage
