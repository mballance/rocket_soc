
`include "uvm_macros.svh"

package rocket_soc_env_pkg;
	import uvm_pkg::*;
	import RocketSocTBEnvBasePkg::*;

	`include "rocket_soc_env.svh"
	
endpackage
